----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Adri�n Hern�ndez
-- Ejercicio 1.19
-- Create Date:    22:30:40 05/23/2022 
-- Design Name: 
-- Module Name:    Robot - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Robot is
    Port ( A,B,C,D : in  STD_LOGIC;
           F : out  STD_LOGIC);
end Robot;

architecture Behavioral of Robot is
begin
	F <= '1' when (A = '1' and B = '1' and C = '1' and D = '1') else '0';

end Behavioral;

